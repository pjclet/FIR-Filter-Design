parameter N_TAPS = 168;