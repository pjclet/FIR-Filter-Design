parameter logic signed[15:0] filter_coeffs[0:167] = '{
16'b1111111111111000,
16'b1111111111101100,
16'b1111111111010000,
16'b1111111110110000,
16'b1111111110000100,
16'b1111111101011100,
16'b1111111100111100,
16'b1111111100110100,
16'b1111111101001000,
16'b1111111101110100,
16'b1111111110111100,
16'b0000000000001000,
16'b0000000001001000,
16'b0000000001101100,
16'b0000000001101100,
16'b0000000001001000,
16'b0000000000001100,
16'b1111111111001100,
16'b1111111110100100,
16'b1111111110100000,
16'b1111111111000000,
16'b1111111111111000,
16'b0000000000111000,
16'b0000000001100000,
16'b0000000001100100,
16'b0000000000111100,
16'b1111111111111100,
16'b1111111110111000,
16'b1111111110010000,
16'b1111111110010100,
16'b1111111111001000,
16'b0000000000010100,
16'b0000000001011100,
16'b0000000010000100,
16'b0000000001110100,
16'b0000000000110100,
16'b1111111111011000,
16'b1111111110000100,
16'b1111111101100000,
16'b1111111110000000,
16'b1111111111011000,
16'b0000000001001000,
16'b0000000010100000,
16'b0000000010111100,
16'b0000000010001100,
16'b0000000000011000,
16'b1111111110010000,
16'b1111111100110000,
16'b1111111100100000,
16'b1111111101110000,
16'b0000000000000100,
16'b0000000010100100,
16'b0000000100001100,
16'b0000000100001000,
16'b0000000010010100,
16'b1111111111010000,
16'b1111111100010100,
16'b1111111010101000,
16'b1111111011001000,
16'b1111111101110100,
16'b0000000001110000,
16'b0000000101010100,
16'b0000000110111100,
16'b0000000101110000,
16'b0000000001110100,
16'b1111111100101000,
16'b1111111000010000,
16'b1111110110110000,
16'b1111111001001000,
16'b1111111110111100,
16'b0000000110001100,
16'b0000001011111000,
16'b0000001101001100,
16'b0000001000110000,
16'b1111111111010000,
16'b1111110011110100,
16'b1111101011000000,
16'b1111101001100100,
16'b1111110010101000,
16'b0000000110101100,
16'b0000100010101100,
16'b0001000000111100,
16'b0001011010100000,
16'b0001101001001000,
16'b0001101001001000,
16'b0001011010100000,
16'b0001000000111100,
16'b0000100010101100,
16'b0000000110101100,
16'b1111110010101000,
16'b1111101001100100,
16'b1111101011000000,
16'b1111110011110100,
16'b1111111111010000,
16'b0000001000110000,
16'b0000001101001100,
16'b0000001011111000,
16'b0000000110001100,
16'b1111111110111100,
16'b1111111001001000,
16'b1111110110110000,
16'b1111111000010000,
16'b1111111100101000,
16'b0000000001110100,
16'b0000000101110000,
16'b0000000110111100,
16'b0000000101010100,
16'b0000000001110000,
16'b1111111101110100,
16'b1111111011001000,
16'b1111111010101000,
16'b1111111100010100,
16'b1111111111010000,
16'b0000000010010100,
16'b0000000100001000,
16'b0000000100001100,
16'b0000000010100100,
16'b0000000000000100,
16'b1111111101110000,
16'b1111111100100000,
16'b1111111100110000,
16'b1111111110010000,
16'b0000000000011000,
16'b0000000010001100,
16'b0000000010111100,
16'b0000000010100000,
16'b0000000001001000,
16'b1111111111011000,
16'b1111111110000000,
16'b1111111101100000,
16'b1111111110000100,
16'b1111111111011000,
16'b0000000000110100,
16'b0000000001110100,
16'b0000000010000100,
16'b0000000001011100,
16'b0000000000010100,
16'b1111111111001000,
16'b1111111110010100,
16'b1111111110010000,
16'b1111111110111000,
16'b1111111111111100,
16'b0000000000111100,
16'b0000000001100100,
16'b0000000001100000,
16'b0000000000111000,
16'b1111111111111000,
16'b1111111111000000,
16'b1111111110100000,
16'b1111111110100100,
16'b1111111111001100,
16'b0000000000001100,
16'b0000000001001000,
16'b0000000001101100,
16'b0000000001101100,
16'b0000000001001000,
16'b0000000000001000,
16'b1111111110111100,
16'b1111111101110100,
16'b1111111101001000,
16'b1111111100110100,
16'b1111111100111100,
16'b1111111101011100,
16'b1111111110000100,
16'b1111111110110000,
16'b1111111111010000,
16'b1111111111101100,
16'b1111111111111000
};
